`timescale 1ns/100ps
`define FAST_SIM
`include "Top.sv"
`include "Random.sv"
`include "DE2_115/SevenHexDecoder.sv"
`include "DE2_115/Debounce.sv"
`include "DE2_115/DE2_115.sv"
