
// CLOCK: 12MHz => 83.33 ns ~= 84 ns
module LCD(
  input        i_clk,
  input        i_rst,
  // LCD module connection
  inout  [7:0] LCD_DATA,
  output       LCD_EN,
  output       LCD_RW,
  output       LCD_RS,
  output       LCD_ON,
  output       LCD_BLON,
  // self designed inout
  output       READY
);

//=======================================================
//-----------------Default Assumption--------------------
//=======================================================

// LCD modules used on DE2-115 boards do not have backlight.
assign LCD_BLON = 1'b0;

//=======================================================
//------------Define Basic Instruction Set---------------
//=======================================================

parameter [7:0] CLEAR      = 8'b00000001; // Execution time = 1.53ms, Clear Display
parameter [7:0] ENTRY_N    = 8'b00000110; // Execution time = 39us,   Normal Entry, Cursor increments, Display is not shifted
parameter [7:0] DISPLAY_ON = 8'b00001100; // Execution time = 39us,   Turn ON Display
parameter [7:0] FUNCT_SET  = 8'b00111000; // Execution time = 39us,   sets to 8-bit interface, 2-line display, 5x8 dots

//=======================================================
//--------------Define Timing Parameters-----------------
//=======================================================

parameter [19:0] t_39us     = 465       //39us      ~= 465    clks
parameter [19:0] t_43us     = 512       //43us      ~= 512    clks
parameter [19:0] t_100us    = 1191;     //100us     ~= 1191   clks
parameter [19:0] t_4100us   = 48810;    //4.1ms     ~= 48810  clks
parameter [19:0] t_15000us  = 178572;   //15ms      ~= 178572 clks

// time counter
logic [19:0] timer_w, timer_r;
logic flag_timer_rst_w, flag_timer_rst_r;
logic flag_39us;
logic flag_43us;
logic flag_100us;
logic flag_4100us;
logic flag_15000us;

//=======================================================
//-------------------Define States-----------------------
//=======================================================

enum {INIT, IDLE, RECORD, STOP, PLAY, PAUSE} state_w, state_r;
enum {SUB_1, SUB_2, SUB_3, SUB_4, SUB_5, SUB_6, SUB_7, SUB_8} substate_w, substate_r;

//=======================================================
//--------------------Time Counter-----------------------
//=======================================================

always_comb begin
  state_w          = state_r;
  substate_w       = substate_r;
  timer_w          = timer_r + 1;
  flag_timer_rst_w = flag_timer_rst_r;
end

always_ff @(posedge i_clk) begin
  if (flag_timer_rst_w) begin
    timer_r      <= 20'b0;
    flag_39us    <= 1'b0;
    flag_43us    <= 1'b0;
    flag_100us   <= 1'b0;
    flag_4100us  <= 1'b0;
    flag_15000us <= 1'b0;
  end else begin
    timer_r <= timer_w;

    if (timer_w >= t_39us) begin
      flag_39us <= 1'b1;
    end else begin
      flag_39us <= flag_39us;
    end

    if (timer_w >= t_43us) begin
      flag_43us <= 1'b1;
    end else begin
      flag_43us <= flag_43us;
    end

    if (timer_w >= t_100us) begin
      flag_100us <= 1'b1;
    end else begin
      flag_100us <= flag_100us;
    end

    if (timer_w >= t_4100us) begin
      flag_4100us <= 1'b1;
    end else begin
      flag_4100us <= flag_4100us;
    end

    if (timer_w >= t_15000us) begin
      flag_15000us <= 1'b1;
    end else begin
      flag_15000us <= flag_15000us;
    end
  end
end


always_ff @(posedge i_clk) begin
  case(state_w)
    INIT: begin
      case(substate_w)
        SUB_1: begin // wait 15ms after Vcc rises to 4.5V
          LCD_DATA <= 8'b0;
          LCD_EN   <= 1'b0;
          LCD_RW   <= 1'b0;
          LCD_RS   <= 1'b0;
          LCD_ON   <= 1'b0;
          READY    <= 1'b0;
          if (!flag_15000us) begin
            substate_r <= substate_w;
            flag_timer_rst_r <= 1'b0;
          end else begin
            substate_r <= SUB_2;
            flag_timer_rst_r <= 1'b1;
          end
        end

        SUB_2: begin // wait for more than 4.1ms
          LCD_DATA <= FUNCT_SET;
          LCD_EN   <= 1'b0;
          LCD_RW   <= 1'b0;
          LCD_RS   <= 1'b0;
          LCD_ON   <= 1'b0;
          READY    <= 1'b0;
        end

        SUB_3: begin
        end

        SUB_4: begin
        end

        SUB_5: begin
        end

        SUB_6: begin
        end

        SUB_7: begin
        end

        SUB_8: begin
        end
    end

    IDLE: begin
    end

    RECORD: begin
    end
    
    STOP: begin
    end
    
    PLAY: begin
    end
    
    PAUSE: begin
    end
end

always_ff @(posedge i_clk or posedge i_rst) begin
  if (i_rst) begin
    state_r        <= INIT;
    substate_r     <= SUB_1;
    flag_timer_rst_r <= 1'b1;
  end
end



endmodule